interface my_if(
    input       clk,
    input       rst_n,
    input [7:0] data,
    input       valid
);

endinterface: my_if
